class moqanitor
endclass
